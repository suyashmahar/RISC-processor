`timescale 1ns / 1ps

module ProcessorTestbench;
   
   reg clk;
   reg RESET;
   reg IRQ;
   
   wire [31:0] InstAdd;
   wire        isCorrect;
   wire [31:0] expAddress;

   integer     i = 0;
   reg [31:0]  ver[1023:0];
   
   assign expAddress = ver[i];
   assign isCorrect = (InstAdd == ver[i]);
      
   Processor uut
     (
      .clk(clk),
      .RESET(RESET),
      .IRQ(IRQ),
      
      .InstAdd(InstAdd)
      );
   
   initial begin
       clk = 1;
       RESET = 0;
       IRQ = 0;
              
       ver[0] = 32'h80000000;
       ver[1] = 32'h8000002C;
       ver[2] = 32'h80000030;
       ver[3] = 32'h80000034;
       ver[4] = 32'h80000038;
       ver[5] = 32'h8000003C;
       ver[6] = 32'h80000040;
       ver[7] = 32'h80000044;
       ver[8] = 32'h80000048;
       ver[9] = 32'h8000004C;
       ver[10] = 32'h80000050;
       ver[11] = 32'h80000054;
       ver[12] = 32'h80000058;
       ver[13] = 32'h8000005C;
       ver[14] = 32'h80000060;
       ver[15] = 32'h80000064;
       ver[16] = 32'h80000068;
       ver[17] = 32'h8000006C;
       ver[18] = 32'h80000070;
       ver[19] = 32'h80000074;
       ver[20] = 32'h80000078;
       ver[21] = 32'h8000007C;
       ver[22] = 32'h80000080;
       ver[23] = 32'h80000084;
       ver[24] = 32'h80000088;
       ver[25] = 32'h8000008C;
       ver[26] = 32'h80000090;
       ver[27] = 32'h80000094;
       ver[28] = 32'h80000098;
       ver[29] = 32'h8000009C;
       ver[30] = 32'h800000A0;
       ver[31] = 32'h800000A4;
       ver[32] = 32'h800000A8;
       ver[33] = 32'h800000AC;
       ver[34] = 32'h800000B0;
       ver[35] = 32'h800000B4;
       ver[36] = 32'h800000B8;
       ver[37] = 32'h800000BC;
       ver[38] = 32'h800000C0;
       ver[39] = 32'h800000C4;
       ver[40] = 32'h800000C8;
       ver[41] = 32'h800000CC;
       ver[42] = 32'h800000D0;
       ver[43] = 32'h800000D4;
       ver[44] = 32'h800000D8;
       ver[45] = 32'h800000DC;
       ver[46] = 32'h800000E0;
       ver[47] = 32'h800000E4;
       ver[48] = 32'h800000E8;
       ver[49] = 32'h800000EC;
       ver[50] = 32'h800000F0;
       ver[51] = 32'h800000F4;
       ver[52] = 32'h800000F8;
       ver[53] = 32'h800000FC;
       ver[54] = 32'h80000100;
       ver[55] = 32'h80000104;
       ver[56] = 32'h80000108;
       ver[57] = 32'h8000010C;
       ver[58] = 32'h80000110;
       ver[59] = 32'h80000114;
       ver[60] = 32'h80000118;
       ver[61] = 32'h8000011C;
       ver[62] = 32'h80000120;
       ver[63] = 32'h80000124;
       ver[64] = 32'h80000128;
       ver[65] = 32'h8000012C;
       ver[66] = 32'h80000130;
       ver[67] = 32'h80000134;
       ver[68] = 32'h80000138;
       ver[69] = 32'h8000013C;
       ver[70] = 32'h80000140;
       ver[71] = 32'h80000144;
       ver[72] = 32'h80000148;
       ver[73] = 32'h8000014C;
       ver[74] = 32'h80000150;
       ver[75] = 32'h80000154;
       ver[76] = 32'h80000158;
       ver[77] = 32'h8000015C;
       ver[78] = 32'h80000160;
       ver[79] = 32'h80000164;
       ver[80] = 32'h80000168;
       ver[81] = 32'h8000016C;
       ver[82] = 32'h80000170;
       ver[83] = 32'h80000174;
       ver[84] = 32'h80000178;
       ver[85] = 32'h8000017C;
       ver[86] = 32'h80000180;
       ver[87] = 32'h80000184;
       ver[88] = 32'h80000188;
       ver[89] = 32'h8000018C;
       ver[90] = 32'h80000190;
       ver[91] = 32'h80000194;
       ver[92] = 32'h80000198;
       ver[93] = 32'h8000019C;
       ver[94] = 32'h800001A0;
       ver[95] = 32'h800001A4;
       ver[96] = 32'h800001A8;
       ver[97] = 32'h800001AC;
       ver[98] = 32'h800001B0;
       ver[99] = 32'h800001B4;
       ver[100] = 32'h800001B8;
       ver[101] = 32'h800001BC;
       ver[102] = 32'h800001C0;
       ver[103] = 32'h800001C4;
       ver[104] = 32'h800001C8;
       ver[105] = 32'h800001CC;
       ver[106] = 32'h800001D0;
       ver[107] = 32'h800001D4;
       ver[108] = 32'h800001D8;
       ver[109] = 32'h800001DC;
       ver[110] = 32'h800001E0;
       ver[111] = 32'h800001E4;
       ver[112] = 32'h800001E8;
       ver[113] = 32'h800001EC;
       ver[114] = 32'h800001F0;
       ver[115] = 32'h800001F4;
       ver[116] = 32'h800001F8;
       ver[117] = 32'h800001FC;
       ver[118] = 32'h80000200;
       ver[119] = 32'h80000204;
       ver[120] = 32'h80000208;
       ver[121] = 32'h8000020C;
       ver[122] = 32'h80000210;
       ver[123] = 32'h80000214;
       ver[124] = 32'h80000218;
       ver[125] = 32'h8000021C;
       ver[126] = 32'h80000220;
       ver[127] = 32'h80000228;
       ver[128] = 32'h8000022C;
       ver[129] = 32'h80000230;
       ver[130] = 32'h80000234;
       ver[131] = 32'h80000238;
       ver[132] = 32'h8000023C;
       ver[133] = 32'h80000240;
       ver[134] = 32'h80000244;
       ver[135] = 32'h80000248;
       ver[136] = 32'h8000024C;
       ver[137] = 32'h80000250;
       ver[138] = 32'h80000254;
       ver[139] = 32'h80000258;
       ver[140] = 32'h8000025C;
       ver[141] = 32'h80000260;
       ver[142] = 32'h80000264;
       ver[143] = 32'h80000268;
       ver[144] = 32'h8000026C;
       ver[145] = 32'h80000270;
       ver[146] = 32'h80000274;
       ver[147] = 32'h80000278;
       ver[148] = 32'h8000027C;
       ver[149] = 32'h80000280;
       ver[150] = 32'h80000284;
       ver[151] = 32'h80000288;
       ver[152] = 32'h8000028C;
       ver[153] = 32'h80000290;
       ver[154] = 32'h80000294;
       ver[155] = 32'h80000298;
       ver[156] = 32'h8000029C;
       ver[157] = 32'h800002A0;
       ver[158] = 32'h800002A4;
       ver[159] = 32'h800002A8;
       ver[160] = 32'h800002AC;
       ver[161] = 32'h800002B0;
       ver[162] = 32'h800002B4;
       ver[163] = 32'h800002B8;
       ver[164] = 32'h800002BC;
       ver[165] = 32'h800002C0;
       ver[166] = 32'h800002C4;
       ver[167] = 32'h800002C8;
       ver[168] = 32'h800002CC;
       ver[169] = 32'h800002D0;
       ver[170] = 32'h800002D4;
       ver[171] = 32'h80000004;
       ver[172] = 32'h80000014;
       ver[173] = 32'h80000018;
       ver[174] = 32'h80000024;
       ver[175] = 32'h80000028;
       ver[176] = 32'h800002D8;
       ver[177] = 32'h800002DC;
       ver[178] = 32'h800002E0;
       ver[179] = 32'h800002E4;
       ver[180] = 32'h800002E8;
       ver[181] = 32'h80000004;
       ver[182] = 32'h80000014;
       ver[183] = 32'h80000018;
       ver[184] = 32'h80000024;
       ver[185] = 32'h80000028;
       ver[186] = 32'h800002EC;
       ver[187] = 32'h80000004;
       ver[188] = 32'h80000014;
       ver[189] = 32'h80000018;
       ver[190] = 32'h80000024;
       ver[191] = 32'h80000028;
       ver[192] = 32'h800002F0;
       ver[193] = 32'h80000004;
       ver[194] = 32'h80000014;
       ver[195] = 32'h80000018;
       ver[196] = 32'h80000024;
       ver[197] = 32'h80000028;
       ver[198] = 32'h800002F4;
       ver[199] = 32'h80000004;
       ver[200] = 32'h80000014;
       ver[201] = 32'h80000018;
       ver[202] = 32'h80000024;
       ver[203] = 32'h80000028;
       ver[204] = 32'h800002F8;
       ver[205] = 32'h80000004;
       ver[206] = 32'h80000014;
       ver[207] = 32'h80000018;
       ver[208] = 32'h80000024;
       ver[209] = 32'h80000028;
       ver[210] = 32'h800002FC;
       ver[211] = 32'h80000004;
       ver[212] = 32'h80000014;
       ver[213] = 32'h80000018;
       ver[214] = 32'h80000024;
       ver[215] = 32'h80000028;
       ver[216] = 32'h80000300;
       ver[217] = 32'h80000004;
       ver[218] = 32'h80000014;
       ver[219] = 32'h80000018;
       ver[220] = 32'h80000024;
       ver[221] = 32'h80000028;
       ver[222] = 32'h80000304;
       ver[223] = 32'h80000004;
       ver[224] = 32'h80000014;
       ver[225] = 32'h80000018;
       ver[226] = 32'h80000024;
       ver[227] = 32'h80000028;
       ver[228] = 32'h80000308;
       ver[229] = 32'h8000030C;
       ver[230] = 32'h80000310;
       ver[231] = 32'h80000314;
       ver[232] = 32'h80000318;
       ver[233] = 32'h8000031C;
       ver[234] = 32'h80000320;
       ver[235] = 32'h80000324;
       ver[236] = 32'h80000328;
       ver[237] = 32'h8000032C;
       ver[238] = 32'h80000330;
       ver[239] = 32'h80000334;
       ver[240] = 32'h80000338;
       ver[241] = 32'h8000033C;
       ver[242] = 32'h80000340;
       ver[243] = 32'h80000344;
       ver[244] = 32'h80000348;
       ver[245] = 32'h8000034C;
       ver[246] = 32'h80000350;
       ver[247] = 32'h80000354;
       ver[248] = 32'h80000358;
       ver[249] = 32'h8000035C;
       ver[250] = 32'h80000360;
       ver[251] = 32'h80000364;
       ver[252] = 32'h80000368;
       ver[253] = 32'h8000036C;
       ver[254] = 32'h80000370;
       ver[255] = 32'h80000374;
       ver[256] = 32'h80000378;
       ver[257] = 32'h8000037C;
       ver[258] = 32'h80000380;
       ver[259] = 32'h80000384;
       ver[260] = 32'h80000388;
       ver[261] = 32'h8000038C;
       ver[262] = 32'h80000390;
       ver[263] = 32'h80000394;
       ver[264] = 32'h80000398;
       ver[265] = 32'h8000039C;
       ver[266] = 32'h800003A0;
       ver[267] = 32'h800003A4;
       ver[268] = 32'h800003A8;
       ver[269] = 32'h800003AC;
       ver[270] = 32'h800003B0;
       ver[271] = 32'h800003B4;
       ver[272] = 32'h000003B8;
       ver[273] = 32'h80000008;
       ver[274] = 32'h000003BC;
       ver[275] = 32'h000003C0;
       ver[276] = 32'h000003C4;
       ver[277] = 32'h000003C8;
       ver[278] = 32'h000003C4;
       ver[279] = 32'h000003C8;
       ver[280] = 32'h000003C4;
       ver[281] = 32'h000003C8;
       ver[282] = 32'h000003C4;
       ver[283] = 32'h000003C8;
       ver[284] = 32'h000003C4;
       ver[285] = 32'h000003C8;
       ver[286] = 32'h000003C4;
       ver[287] = 32'h000003C8;     

      #20
	RESET = 1;
      #10
	RESET = 0;
   end

   always begin
       #40 clk = ~clk;
   end

   always begin
       #80 
       i = i+1;
   end

   always begin
       #21820
	 IRQ = ~IRQ;
       #25 
	 IRQ = ~IRQ;
   end

   

   always begin
       #2000
	 IRQ = ~IRQ;
       #100
	 IRQ = ~IRQ;
   end
endmodule // ProcessorTestbench

