`timescale 1ns / 1ps

module Shifter_Testbench;

reg [5:0] alufn;
reg [31:0] a;
reg [31:0] b;

wire [31:0] s;
wire z;
wire v;
wire n;

wire [31:0] shtRes;
reg [31:0] isCorrect;
reg [31:0] expRes;



reg [99:0] val [95:0];

integer i = 0;

ShifterModule shft_inst_0 (
    .alufn(alufn),
    .a(a),
    .b(b),

    .res(shtRes)
);

initial begin 
    //            <-res--> <--a---> <--b---> allufn[4:0]
    val[0] = 100'h87654321_87654321_00000000_0;
    val[1] = 100'h0ECA8642_87654321_00000001_0;
    val[2] = 100'h1D950C84_87654321_00000002_0;
    val[3] = 100'h3B2A1908_87654321_00000003_0;
    val[4] = 100'h76543210_87654321_00000004_0;
    val[5] = 100'hECA86420_87654321_00000005_0;
    val[6] = 100'hD950C840_87654321_00000006_0;
    val[7] = 100'hB2A19080_87654321_00000007_0;
    val[8] = 100'h65432100_87654321_00000008_0;
    val[9] = 100'hCA864200_87654321_00000009_0;
    val[10] = 100'h950C8400_87654321_0000000A_0;
    val[11] = 100'h2A190800_87654321_0000000B_0;
    val[12] = 100'h54321000_87654321_0000000C_0;
    val[13] = 100'hA8642000_87654321_0000000D_0;
    val[14] = 100'h50C84000_87654321_0000000E_0;
    val[15] = 100'hA1908000_87654321_0000000F_0;
    val[16] = 100'h43210000_87654321_00000010_0;
    val[17] = 100'h86420000_87654321_00000011_0;
    val[18] = 100'h0C840000_87654321_00000012_0;
    val[19] = 100'h19080000_87654321_00000013_0;
    val[20] = 100'h32100000_87654321_00000014_0;
    val[21] = 100'h64200000_87654321_00000015_0;
    val[22] = 100'hC8400000_87654321_00000016_0;
    val[23] = 100'h90800000_87654321_00000017_0;
    val[24] = 100'h21000000_87654321_00000018_0;
    val[25] = 100'h42000000_87654321_00000019_0;
    val[26] = 100'h84000000_87654321_0000001A_0;
    val[27] = 100'h08000000_87654321_0000001B_0;
    val[28] = 100'h10000000_87654321_0000001C_0;
    val[29] = 100'h20000000_87654321_0000001D_0;
    val[30] = 100'h40000000_87654321_0000001E_0;
    val[31] = 100'h80000000_87654321_0000001F_0;
    val[32] = 100'hFEDCBA98_FEDCBA98_00000000_1;
    val[33] = 100'h3F6E5D4C_7EDCBA98_00000001_1;
    val[34] = 100'h3FB72EA6_FEDCBA98_00000002_1;
    val[35] = 100'h0FDB9753_7EDCBA98_00000003_1;
    val[36] = 100'h0FEDCBA9_FEDCBA98_00000004_1;
    val[37] = 100'h03F6E5D4_7EDCBA98_00000005_1;
    val[38] = 100'h03FB72EA_FEDCBA98_00000006_1;
    val[39] = 100'h00FDB975_7EDCBA98_00000007_1;
    val[40] = 100'h007EDCBA_7EDCBA98_00000008_1;
    val[41] = 100'h007F6E5D_FEDCBA98_00000009_1;
    val[42] = 100'h001FB72E_7EDCBA98_0000000A_1;
    val[43] = 100'h001FDB97_FEDCBA98_0000000B_1;
    val[44] = 100'h0007EDCB_7EDCBA98_0000000C_1;
    val[45] = 100'h0007F6E5_FEDCBA98_0000000D_1;
    val[46] = 100'h0001FB72_7EDCBA98_0000000E_1;
    val[47] = 100'h0001FDB9_FEDCBA98_0000000F_1;
    val[48] = 100'h0000FEDC_FEDCBA98_00000010_1;
    val[49] = 100'h00003F6E_7EDCBA98_00000011_1;
    val[50] = 100'h00003FB7_FEDCBA98_00000012_1;
    val[51] = 100'h00000FDB_7EDCBA98_00000013_1;
    val[52] = 100'h00000FED_FEDCBA98_00000014_1;
    val[53] = 100'h000003F6_7EDCBA98_00000015_1;
    val[54] = 100'h000003FB_FEDCBA98_00000016_1;
    val[55] = 100'h000000FD_7EDCBA98_00000017_1;
    val[56] = 100'h0000007E_7EDCBA98_00000018_1;
    val[57] = 100'h0000007F_FEDCBA98_00000019_1;
    val[58] = 100'h0000001F_7EDCBA98_0000001A_1;
    val[59] = 100'h0000001F_FEDCBA98_0000001B_1;
    val[60] = 100'h00000007_7EDCBA98_0000001C_1;
    val[61] = 100'h00000007_FEDCBA98_0000001D_1;
    val[62] = 100'h00000001_7EDCBA98_0000001E_1;
    val[63] = 100'h00000001_FEDCBA98_0000001F_1;
    val[64] = 100'h87654321_87654321_00000000_3;
    val[65] = 100'h3B2A1908_76543210_00000001_3;
    val[66] = 100'hE1D950C8_87654321_00000002_3;
    val[67] = 100'h0ECA8642_76543210_00000003_3;
    val[68] = 100'hF8765432_87654321_00000004_3;
    val[69] = 100'h03B2A190_76543210_00000005_3;
    val[70] = 100'hFE1D950C_87654321_00000006_3;
    val[71] = 100'h00ECA864_76543210_00000007_3;
    val[72] = 100'h00765432_76543210_00000008_3;
    val[73] = 100'hFFC3B2A1_87654321_00000009_3;
    val[74] = 100'h001D950C_76543210_0000000A_3;
    val[75] = 100'hFFF0ECA8_87654321_0000000B_3;
    val[76] = 100'h00076543_76543210_0000000C_3;
    val[77] = 100'hFFFC3B2A_87654321_0000000D_3;
    val[78] = 100'h0001D950_76543210_0000000E_3;
    val[79] = 100'hFFFF0ECA_87654321_0000000F_3;
    val[80] = 100'hFFFF8765_87654321_00000010_3;
    val[81] = 100'h00003B2A_76543210_00000011_3;
    val[82] = 100'hFFFFE1D9_87654321_00000012_3;
    val[83] = 100'h00000ECA_76543210_00000013_3;
    val[84] = 100'hFFFFF876_87654321_00000014_3;
    val[85] = 100'h000003B2_76543210_00000015_3;
    val[86] = 100'hFFFFFE1D_87654321_00000016_3;
    val[87] = 100'h000000EC_76543210_00000017_3;
    val[88] = 100'h00000076_76543210_00000018_3;
    val[89] = 100'hFFFFFFC3_87654321_00000019_3;
    val[90] = 100'h0000001D_76543210_0000001A_3;
    val[91] = 100'hFFFFFFF0_87654321_0000001B_3;
    val[92] = 100'h00000007_76543210_0000001C_3;
    val[93] = 100'hFFFFFFFC_87654321_0000001D_3;
    val[94] = 100'h00000001_76543210_0000001E_3;
    val[95] = 100'hFFFFFFFF_87654321_0000001F_3;
end

always begin
    #10
    i = i + 1;
    alufn = {{3'b0}, {val[i][1:0]}};
    a = val[i][67:36];
    b = val[i][35:4];
    expRes = val[i][99:68];
    isCorrect = ~(shtRes == val[i][99:68]);
end
endmodule
